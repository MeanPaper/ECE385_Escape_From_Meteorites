module random_generater(input[9:0] randomX, randomY,	//random x and y position
								input[3:0] random_x_speed, random_y_speed,	//random x and y speed
								input object_alive[4],	//activation record
								output[9:0] new_obj_x[4], new_obj_y[4],	//new position of the objects
								output[3:0] new_x_speed[4], new_y_speed[4]	//new speed of the objects
								);
								


endmodule
