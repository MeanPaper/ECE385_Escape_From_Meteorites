module counter_rand(input Clk);

endmodule
